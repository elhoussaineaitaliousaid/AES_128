library ieee;
use ieee.std_logic_1164.all;

package types_pkg is
    type array_bytes is array(0 to 15) of std_logic_vector(7 downto 0);
end package;

package body types_pkg is
end package body;
